/* Definition of the `ping` component. */

component forte.NavigationCommand

endpoints {
    /* Declaration of a named implementation of the "Ping" interface. */
    setNavigationCommand : forte.NavigationCommand
}
